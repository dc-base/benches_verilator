`include "full_adder.sv"
`include "barrel_shifter.sv"
`include "multiplier.sv"

module alu_control()


endmodule
